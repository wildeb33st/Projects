library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.coeff_pkg.all; 

entity test_bench is
--  Port ( );
end test_bench;



architecture a of test_bench is
-- VALIDATE THESE CLOCK TIMES!!!!!!!
    constant CLOCK_PERIOD    : time := 50  ps;
    constant SIMULATION_TIME : time := 1000 ps;

    signal clk      : std_logic := '0';
    
---------------------------------------------------------------------------------------------------------------------------------
--Below are interconnecting signals etc. for components

-- This is for the read line for taking data from fileRd component output (data)
-- to DUT component input (din)
    signal readLn :  integer := 0;
    
--signal for reading imaginary components from file    
    signal readLnIm : integer := 0;
    
--Write line signal is used for moving data from the output of the DUT component
-- to the input of the fileWr component
    signal writeLn : integer := 0;

--input to the file for Imaginary Filter output    
    signal writeLnIm : integer := 0;

--DV line for the purpose of letting DUT know when a signal is incoming
    signal dvLn : std_logic := '1';

-- Reset signal for reader
signal rst    : std_logic := '0';

--Rfd signal for reader
signal rfd : std_logic := '1';

--constant for reader to state bit width
constant numOfBits : integer := 16;

--constant for readfile
constant file_name : string := "/home/gear/Downloads/ProjectFilter/data2fpga2.dat";

--constant for readfile Imaginary Filter
constant file_nameIm : string := "/home/gear/Downloads/ProjectFilter/data2fpga_imag.dat";

--constant for written file
constant file_name_wr : string := "/home/gear/Downloads/ProjectFilter/data_from_fpga.dat";

--constant for written file
constant file_name_wrIm : string := "/home/gear/Downloads/ProjectFilter/data_from_fpga_Im.dat";

--Constants for the filter are below
constant input_width :integer:=16;-- this is based on the input data width 
constant output_width:integer:=32;-- this is twice the size since the coefficient will be the same size
constant coef_width:integer:=16;--Barker code is used as coefficient and is converted to 16-bit width
constant tap:integer:=13; --11-chip barker sequence was specified and so this is used

--constant representing the coefficient for the real filter
constant coeficient : Coeficient_type := (1, -1, 1, -1, 1, 1, -1, -1, 1, 1, 1, 1, 1);

----constant representing the coefficient for the Imaginary filter
constant coeficientIm : Coeficient_type := (-1, 1, -1, 1, -1, -1, 1, 1, -1, -1, -1, -1, -1);

----------------------------------------------------------------------------------------------------------------------------------
--Components

--Lab12 Component i.e. The Device Under Test (DUT)
    component FIR_RI is
        generic (  
--           input_width :integer:=16;-- this is based on the input data width 
--           output_width:integer:=32;-- this is twice the size since the coefficient will be the same size
--           coef_width:integer:=16;--Barker code is used as coefficient and is converted to 16-bit width
           tap:integer:=11; --11-chip barker sequence was specified and so this is used
           coeficient : Coeficient_type
         );    
        port(
            Din:in integer; -- input data 
            Clk:in std_logic; -- input clk  
            reset:in std_logic; -- input reset  
            Dout:out integer -- output data
            );
    end component FIR_RI;

--Component to read the Sine Wave Amplitude Values that were generated by MATLAB Script
component ReadFile is
        generic(
         --        numOfBits : integer;
                 file_name : string
               );
        Port (
                data : out integer;
                dv: out std_logic;
                rst : in std_logic;
                rfd : in std_logic;
                clk : in std_logic
              );
end component ReadFile;

--Component for writing FPGA results to another file
component WriteFile_full
        generic(
                 --output_width : integer;
                 file_name : string
               );
        Port (
                clk,dv : in std_logic;
                DataIn : in integer
              );
end component WriteFile_full;

----------------------------------------------------------------------------------------------------------------------------------------

begin

  -----------------------------------------------------------------------
  -- Generate clock
  -----------------------------------------------------------------------
  clock_gen : process
  begin
    clk <= '0';
    wait for CLOCK_PERIOD;
    loop
      clk <= '1';
      wait for CLOCK_PERIOD/2;
      clk <= '0';
      wait for CLOCK_PERIOD/2;
    end loop;
  end process clock_gen;
  -----------------------------------------------------------------------
  -- Generate start
  -----------------------------------------------------------------------
  start_gen : process
  begin
    rst <= '1';
    wait for CLOCK_PERIOD;
    wait for CLOCK_PERIOD;
    wait for CLOCK_PERIOD;
    rst <= '0';

    wait for CLOCK_PERIOD;
    rst <= '0';
    wait;
  end process start_gen;

  ---------------------------------------------------------------------
  -- Instantiate the DUT
  ---------------------------------------------------------------------
--  DUT : lab111
--    port map (
--        -- Inputs
--        clk => clk,
--        din => readLn,
--        dv => dvLn,
--        -- Outputs
--        dout  => writeLn);
        
  ---------------------------------------------------------------------
  --Real Filter
  ---------------------------------------------------------------------  
  RealFilter : FIR_RI
     generic map (  
                 --   input_width => input_width, 
                 --   output_width => output_width,
                 --   coef_width => coef_width,
                    tap => tap,
                    coeficient => coeficient
                 )
                     
     port map (
        
              Din => readLn,  
              Clk => clk, 
              reset => rst,  
              Dout => writeLn
            
            );
    


---------------------------------------------------------------------
  --Imaginary Filter
  ---------------------------------------------------------------------  
  ImaginaryFilter : FIR_RI
     generic map (  
                 --   input_width => input_width, 
                 --   output_width => output_width,
                 --   coef_width => coef_width,
                    tap => tap,
                    coeficient => coeficientIm
                 )
                     
     port map (
        
              Din => readLnIm,  
              Clk => clk, 
              reset => rst,  
              Dout => writeLnIm
            
            );
    


  ---------------------------------------------------------------------
  -- Instantiate the Reader to read from file
  ---------------------------------------------------------------------
  reader : ReadFile
    generic map (
                   -- numOfBits => numOfBits,
                    file_name => file_name
                )
    port map (
                data => readLn,
                dv => dvLn,
                clk => clk,
                rst => rst,
                rfd => rfd
              );
              

 ---------------------------------------------------------------------
  -- Instantiate the Reader to read from file (Imaginary Component)
  ---------------------------------------------------------------------
  readerIm : ReadFile
    generic map (
                   -- numOfBits => numOfBits,
                    file_name => file_nameIm
                )
    port map (
                data => readLnIm,
                dv => dvLn,
                clk => clk,
                rst => rst,
                rfd => rfd
              );
 

  ---------------------------------------------------------------------
  -- Instantiate the writer to write to a file
  ---------------------------------------------------------------------
  writer : WriteFile_full
    generic map (
                   -- output_width => output_width,
                    file_name => file_name_wr
                )
    port map (
                dv => dvLn,
                clk => clk,
               -- sign => writeLn(31),
                DataIn => writeLn
              );



  ---------------------------------------------------------------------
  -- Instantiate the writer to write to a file
  ---------------------------------------------------------------------
  writerIm : WriteFile_full
    generic map (
                   -- output_width => output_width,
                    file_name => file_name_wrIm
                )
    port map (
                dv => dvLn,
                clk => clk,
               -- sign => writeLn(31),
                DataIn => writeLnIm
              );




end architecture;
                  
